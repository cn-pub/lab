`timescale 1ns / 1ps
module cla_subtractor (
        output  [7: 0] D,
        output                      Cout,
        input   [7: 0] A,
        input   [7: 0] B,
        input                       Cin
    );

    //TODO 2: implemetati logica pentru un scazator carry-lookahead pe 4 biti
endmodule

