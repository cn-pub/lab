// Copyright 2018 Darius Neatu <neatudarius@gmail.com>

`include "defines.vh"

module test_ual;
  `include "tester.vh"

	// outputs
	wire [7:0] out;
	reg  [7:0] expected;

	// Inputs
	reg [4:0] opcode;
	reg [3:0] A;
	reg [3:0] B;

	// spartan stuff
	reg button;
	reg reset;
	reg clk;
	
	// checker
	reg [7:0] respect;
	reg  result;


	reg [1024 * 8 - 1 : 0] opname;

	// Instantiate the Unit Under Test (UUT)
	ual #(.DATA_WIDTH(4) ) uut (
    	.out(out),
		.sel(opcode),
		.in0(A), 
		.in1(B)
	);
	
	initial begin
		clk  = 0;
		
		// Initialize Inputs
		opcode = 0;
		A = 0;
		B = 0;
		
		button = 0;
		reset = 1;
		respect = 0;

		#10;
		reset = 0;
		
		// =======================================================
		// =======================================================
		// TEST NAND: A = 0, B = 0
		#10;
		opname = "NAND";
		opcode = 5'd1;
                  A = 4'b0000;
		            B = 4'b0000;
		expected = 8'b0000_1111;
		#10; 
		if (1'b1 == tester(opname, opcode, expected, out, A, B)) begin
			respect = respect + 1;
		end
		// =======================================================
		// =======================================================
		
		
		// =======================================================
		// =======================================================
		// TEST NAND: A = 15, B = 15
		#10;
		opname = "NAND";
		opcode = 5'd1;
                  A = 4'b1111;
		            B = 4'b1111;
		expected = 8'b0000_0000;
		#10; 
		if (1'b1 == tester(opname, opcode, expected, out, A, B)) begin
			respect = respect + 1;
		end
		// =======================================================
		// =======================================================
		
		
		// =======================================================
		// =======================================================
		// TEST NAND: A = 6, B = 9
		#10;
		opname = "NAND";
		opcode = 5'd1;
                  A = 4'b0110;
		            B = 4'b1001;
		expected = 8'b0000_1111;
		#10; 
		if (1'b1 == tester(opname, opcode, expected, out, A, B)) begin
			respect = respect + 1;
		end
		// =======================================================
		// =======================================================
		
		
		// =======================================================
		// =======================================================
		// TEST XOR: A = 0, B = 0
		#10;
		opname = "XOR";
		opcode = 5'd2;
                  A = 4'b0000;
		            B = 4'b0000;
		expected = 8'b0000_0000;
		#10; 
		if (1'b1 == tester(opname, opcode, expected, out, A, B)) begin
			respect = respect + 1;
		end
		// =======================================================
		// =======================================================
		
		
		// =======================================================
		// =======================================================
		// TEST XOR: A = 3, B = 7
		#10;
		opname = "XOR";
		opcode = 5'd2;
                  A = 4'b0011;
		            B = 4'b0111;
		expected = 8'b0000_0100;
		#10; 
		if (1'b1 == tester(opname, opcode, expected, out, A, B)) begin
			respect = respect + 1;
		end
		// =======================================================
		// =======================================================
		
		
		// =======================================================
		// =======================================================
		// TEST XOR: A = 10, B = 5
		#10;
		opname = "XOR";
		opcode = 5'd2;
                  A = 4'b1010;
		            B = 4'b0101;
		expected = 8'b0000_1111;
		#10; 
		if (1'b1 == tester(opname, opcode, expected, out, A, B)) begin
			respect = respect + 1;
		end
		// =======================================================
		// =======================================================
		
		
		// =======================================================
		// =======================================================
		// TEST ADD: A = 0, B = 0
		#10;
		opname = "ADD";
		opcode = 5'd4;
                  A = 4'b0000;
		            B = 4'b0000;
		expected = 8'b0000_0000;
		#10; 
		if (1'b1 == tester(opname, opcode, expected, out, A, B)) begin
			respect = respect + 1;
		end
		// =======================================================
		// =======================================================
		
		
		
		// =======================================================
		// =======================================================
		// TEST ADD: A = 1, B = 5
		#10;
		opname = "ADD";
		opcode = 5'd4;
                  A = 4'b0001;
		            B = 4'b0101;
		expected = 8'b0000_0110;
		#10; 
		if (1'b1 == tester(opname, opcode, expected, out, A, B)) begin
			respect = respect + 1;
		end
		// =======================================================
		// =======================================================
		
		
		
		// =======================================================
		// =======================================================
		// TEST ADD: A = 5, B = 1
		#10;
		opname = "ADD";
		opcode = 5'd4;
                  A = 4'b0101;
		            B = 4'b0001;
		expected = 8'b0000_0110;
		#10; 
		if (1'b1 == tester(opname, opcode, expected, out, A, B)) begin
			respect = respect + 1;
		end
		// =======================================================
		// =======================================================
		
		
		
		// =======================================================
		// =======================================================
		// TEST ADD: A = 6, B = 9
		#10;
		opname = "ADD";
		opcode = 5'd4;
                  A = 4'b0110;
		            B = 4'b1001;
		expected = 8'b0000_1111;
		#10; 
		if (1'b1 == tester(opname, opcode, expected, out, A, B)) begin
			respect = respect + 1;
		end
		// =======================================================
		// =======================================================
		
		
		// =======================================================
		// =======================================================
		// TEST ADD: A = 6, B = 6
		#10;
		opname = "ADD";
		opcode = 5'd4;
                  A = 4'b0110;
		            B = 4'b0110;
		expected = 8'b0000_1100;
		#10; 
		if (1'b1 == tester(opname, opcode, expected, out, A, B)) begin
			respect = respect + 1;
		end
		// =======================================================
		// =======================================================
		
		
		
		// =======================================================
		// =======================================================
		// TEST SUB: A = 0, B = 0
		#10;
		opname = "SUB";
		opcode = 5'd8;
                  A = 4'b0000;
		            B = 4'b0000;
		expected = 8'b0000_0000;
		#10; 
		if (1'b1 == tester(opname, opcode, expected, out, A, B)) begin
			respect = respect + 1;
		end
		// =======================================================
		// =======================================================
		
		
		
		// =======================================================
		// =======================================================
		// TEST SUB: A = 7, B = 5
		#10;
		opname = "SUB";
		opcode = 5'd8;
                  A = 4'b0111;
		            B = 4'b0101;
		expected = 8'b0000_0010;
		#10; 
		if (1'b1 == tester(opname, opcode, expected, out, A, B)) begin
			respect = respect + 1;
		end
		// =======================================================
		// =======================================================
		
		
		// =======================================================
		// =======================================================
		// TEST SUB: A = 5, B = 7
		#10;
		opname = "SUB";
		opcode = 5'd8;
                  A = 4'b0101;
		            B = 4'b0111;
		expected = 8'b0000_1110;
		#10; 
		if (1'b1 == tester(opname, opcode, expected, out, A, B)) begin
			respect = respect + 1;
		end
		// =======================================================
		// =======================================================
		
		
		// =======================================================
		// =======================================================
		// TEST SUB: A = 2, B = -2
		#10;
		opname = "SUB";
		opcode = 5'd8;
                  A = 4'b0010;
		            B = 4'b1110;
		expected = 8'b0000_0100;
		#10; 
		if (1'b1 == tester(opname, opcode, expected, out, A, B)) begin
			respect = respect + 1;
		end
		// =======================================================
		// =======================================================
		
		
		
		
		// =======================================================
		// =======================================================
		// TEST SUB: A = -2, B = -1
		#10;
		opname = "SUB";
		opcode = 5'd8;
                  A = 4'b1110;
		            B = 4'b1111;
		expected = 8'b0000_1111;
		#10; 
		if (1'b1 == tester(opname, opcode, expected, out, A, B)) begin
			respect = respect + 1;
		end
		// =======================================================
		// =======================================================
		
		

		// =======================================================
		// =======================================================
		// TEST MUL: A = 2, B = 0
		#10;
		opname = "MUL";
		opcode = 5'd16;
             A =      4'b0010;
		       B =      4'b0000;
		expected = 8'b0000_0000;
		#10; 
		if (1'b1 == tester(opname, opcode, expected, out, A, B)) begin
			respect = respect + 1;
		end
		// =======================================================
		// =======================================================
		
		
		
		// =======================================================
		// TEST MUL: A = 2, B = 1
		#10;
		opname = "MUL";
		opcode = 5'd16;
             A =      4'b0010;
		       B =      4'b0001;
		expected = 8'b0000_0010;
		#10; 
		if (1'b1 == tester(opname, opcode, expected, out, A, B)) begin
			respect = respect + 1;
		end
		// =======================================================
		// =======================================================
		
		
		
		// =======================================================
		// TEST MUL: A = 2, B = -1
		#10;
		opname = "MUL";
		opcode = 5'd16;
             A =      4'b0010;
		       B =      4'b1111;
		expected = 8'b1111_1110;
		#10; 
		if (1'b1 == tester(opname, opcode, expected, out, A, B)) begin
			respect = respect + 1;
		end
		// =======================================================
		// =======================================================
		
		
		
		// =======================================================
		// TEST MUL: A = 4, B = 4
		#10;
		opname = "MUL";
		opcode = 5'd16;
             A =      4'b0100;
		       B =      4'b0100;
		expected = 8'b0001_0000;
		#10; 
		if (1'b1 == tester(opname, opcode, expected, out, A, B)) begin
			respect = respect + 1;
		end
		// =======================================================
		// =======================================================
		
		
		
		// =======================================================
		// TEST MUL: A = 4, B = -4
		#10;
		opname = "MUL";
		opcode = 5'd16;
             A =      4'b0100;
		       B =      4'b1100;
		expected = 8'b1111_0000;
		#10; 
		if (1'b1 == tester(opname, opcode, expected, out, A, B)) begin
			respect = respect + 1;
		end
		// =======================================================
		// =======================================================
		
		
		
		// =======================================================
		// TEST MUL: A = -4, B = 4
		#10;
		opname = "MUL";
		opcode = 5'd16;
             A =      4'b1100;
		       B =      4'b0100;
		expected = 8'b1111_0000;
		#10; 
		if (1'b1 == tester(opname, opcode, expected, out, A, B)) begin
			respect = respect + 1;
		end
		// =======================================================
		// =======================================================
		
		
		
		// =======================================================
		// TEST MUL: A = -4, B = -4
		#10;
		opname = "MUL";
		opcode = 5'd16;
             A =      4'b1100;
		       B =      4'b1100;
		expected = 8'b0001_0000;
		#10; 
		if (1'b1 == tester(opname, opcode, expected, out, A, B)) begin
			respect = respect + 1;
		end
		// =======================================================
		// =======================================================
		
		$display("Teste UAL = %2d/23", respect); 
	end
	
	always #1 clk = ~clk;
      
endmodule

