`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    19:44:19 04/05/2020 
// Design Name: 
// Module Name:    adder_32b 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module adder_32b(
    output[31:0] S,
    output Cout,
    input[31:0] A,
    input[31:0] B,
    input Cin
    );

	// TODO 3: Implementati un adder pe 32 de biti (Hint: don't write too much code)
	
endmodule
