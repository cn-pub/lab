`timescale 1ns / 1ps

//////////////////////////////////////////////////////////////////////////////////
// ACS
// Computer Design 1
//  
// Module Name:  		ripple_carry_8bit
// Project Name:		Laborator 6
// Target Devices: 		Digilent Nexys 3
//////////////////////////////////////////////////////////////////////////////////

module ripple_carry_8bit(
		output carry_out,
		output [7:0] sum,
		input  [7:0] A,
		input  [7:0] B,
		input carry_in
    );
	
	// TODO 2: Implementati un sumator ripple-carry pe 8 biti folosind modul full-adder implementat anterior.
	// Hint: buffer pentru transportul din rangul inferior
	
endmodule
