`timescale 1ns / 1ps

//////////////////////////////////////////////////////////////////////////////////
// ACS
// Computer Design 1
//  
// Module Name:  		subtractor_8bit
// Project Name:		Laborator 6
// Target Devices: 		Digilent Nexys 3
//////////////////////////////////////////////////////////////////////////////////

module subtractor_8bit(
		output carry_out,
		output [7:0] result,
		input  [7:0] A,
		input  [7:0] B,
		input carry_in
    );

	// TODO 3: Implementati un sc�z�tor pe 8 biti folosind sumatorul ripple-carry implementat
	// Conventie: result = A - B
	// Hint: Complement fat� de 2
	
endmodule
