module exemplu(
    output out,
    input in
    );

    not(out, in);
	
endmodule
