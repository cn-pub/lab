`timescale 1ns / 1ps

//////////////////////////////////////////////////////////////////////////////////
// ACS
// Computer Design 1
//  
// Module Name:  		full_adder
// Project Name:		Laborator 6
// Target Devices: 		Digilent Nexys 3
//////////////////////////////////////////////////////////////////////////////////

module full_adder(
		output sum,
		output carry_out,
		input bit_A,
		input bit_B,
		input carry_in
    );
	
	// TODO 1.4: Implementati un full-adder folosind dou� instante ale modulului half-adder creat anterior.

endmodule
