`define ZF 4
`define CF 5
`define OF 6
`define SF 7
