module hello_world(
    output led,
    input button
    );

    assign led = button;
endmodule
