// CN1 -  schelet lab02

module modul01(
  output out,
  input in
  );

  not(out, in);

endmodule