/* Constants */
`define SMPHR_RED_TMR				8'd40
`define SMPHR_GRN_TMR				8'd20
`define SMPHR_TMR_START				8'd1
`define SMPHR_TMR_STOP				8'd1
`define OUT_SYNC					8'd1
`define LED_TMR						8'd10

/* Checker */
`define CLK_PERIOD					2
`define EX1_TOTAL					8'd3
`define EX1_SCORE					1.5
`define EX2_TOTAL					8'd17
`define EX2_SCORE					3
`define EX3_TOTAL					8'd4
`define EX3_SCORE					3.5
`define EX4_TOTAL					8'd6
`define EX4_SCORE					4