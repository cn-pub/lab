`timescale 1ns / 1ps
module cla_adder (
        output  [7: 0] S,
        output         Cout,
        input   [7: 0] A,
        input   [7: 0] B,
        input          Cin
    );

	//TODO 1: implemetati logica unui sumator carry-lookahead pe 4 biti,

    
endmodule

